// RISC-V SiMPLE SV -- configuration for testbench
// BSD 3-Clause License
// (c) 2017-2020, Arthur Matos, Marcus Vinicius Lamar, Universidade de Brasília,
//                Marek Materzok, Jakub Piecuch, University of Wrocław

`ifndef RV_CONFIG
`define RV_CONFIG

// Select architecture
`define SINGLE_CYCLE
// `define MULTI_CYCLE
// `define PIPELINE

`include "../common_config.sv"

`endif
